library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity RIGHT_SHIFT_MULTIPLIER is
	generic (
			SIZE : integer := 8  -- Size of the operands
		);
	port (
		     CLOCK     : in  STD_LOGIC;
		     RESET     : in  STD_LOGIC;
		     START     : in  STD_LOGIC;
		     A         : in  STD_LOGIC_VECTOR(SIZE-1 downto 0);
		     B         : in  STD_LOGIC_VECTOR(SIZE-1 downto 0);
		     PRODUCT   : out STD_LOGIC_VECTOR((2*SIZE)-1 downto 0);
		     DONE      : out STD_LOGIC
	     );
end entity;

architecture ARCH of RIGHT_SHIFT_MULTIPLIER is
	signal STATE           : STD_LOGIC_VECTOR(2 downto 0);
	signal NEXT_STATE      : STD_LOGIC_VECTOR(2 downto 0);
	signal MULTIPLICAND    : STD_LOGIC_VECTOR(SIZE-1 downto 0);
	signal PARTIAL_PRODUCT : STD_LOGIC_VECTOR((2*SIZE) downto 0);
	signal ACTIVE          : STD_LOGIC := '0';
	signal ADDER_IN        : STD_LOGIC_VECTOR((2*SIZE)-1 downto 0);
	signal ADDER_OUT       : STD_LOGIC_VECTOR((2*SIZE) downto 0);
begin
	process(CLOCK, RESET)
	begin
		if RESET = '1' then
			MULTIPLICAND    <= (others => '0');
			PARTIAL_PRODUCT <= (others => '0');
			SHIFT_REG       <= (others => '0');
			ACTIVE          <= '0';
		elsif rising_edge(CLOCK) then
			if START = '1' and ACTIVE = '0' then
				MULTIPLICAND    <= B;
				PARTIAL_PRODUCT <= (others => '0');
				PARTIAL_PRODUCT(SIZE-1 downto 0) <= A;
				SHIFT_REG       <= (others => '0');
				ACTIVE          <= '1';
			elsif ACTIVE = '1' then
				if PARTIAL_PRODUCT(1) = '1' then
					ADDER_IN <= MULTIPLICAND & (others => '0');
				else
					ADDER_IN <= (other => '0');
				end if;
				ADDER_OUT <= std_logic_vector(unsigned(PARTIAL_PRODUCT) + unsigned(ADDER_IN));
				PARTIAL_PRODUCT <= ADDER_OUT srl 1;

				case STATE is
					when "000" => NEXT_STATE <= "001";
					when "001" => NEXT_STATE <= "010";
					when "010" => NEXT_STATE <= "011";
					when "011" => NEXT_STATE <= "100";
					when "100" => NEXT_STATE <= "101";
					when "101" => NEXT_STATE <= "110";
					when "110" => NEXT_STATE <= "111";
					when "111" => 
						NEXT_STATE <= "000";
						ACTIVE <= '0';
				end case;
			end if;
		end if;
	end process;

	STATE   <= NEXT_STATE;
	PRODUCT <= PARTIAL_PRODUCT((2*SIZE)-1 downto 0);
	DONE    <= not ACTIVE;

end architecture;
